module decoder_manch #(
    parameter 
) (
  input  wire clk,
  input  wire rx_data,
  output wire tx_data

);
  
  always @(posedge clk) begin
    
  end
    
endmodule